module top (input clk, reset,output [15:0] writedata, dataadr,output memwrite);
wire [15:0] pc, instr, readdata;
// instantiate processor and memories
mips mips (clk, reset, pc, instr, memwrite, dataadr,
writedata, readdata);
imem imem (pc[3:1], instr);
dmem dmem (clk, memwrite, dataadr, writedata,readdata);
endmodule
module branchType (input branch, output btype);
assign btype = branch;
endmodule